`timescale 1ns/100ps

module top_tb();

endmodule
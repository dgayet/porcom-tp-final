module ffe
#(
    parameter NB = 10
)
(
    input i_clock,
    input i_reset
);

endmodule;